module mymodule

// To export a function we have to use `pub`
pub fn hello(name string) string {
	return 'hello $name'
}