// mymodule/mymodule_test.v
module mymodule

fn test_hello() {
	assert hello('tkm') == 'hello tkm'
}